library verilog;
use verilog.vl_types.all;
entity nios_old_tb is
end nios_old_tb;
