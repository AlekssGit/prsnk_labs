library verilog;
use verilog.vl_types.all;
entity nios_old_nios2_qsys_0_nios2_performance_monitors is
end nios_old_nios2_qsys_0_nios2_performance_monitors;
