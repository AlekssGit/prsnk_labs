
module nios (
	board_led_export,
	clk_clk,
	reset_reset_n);	

	output	[3:0]	board_led_export;
	input		clk_clk;
	input		reset_reset_n;
endmodule
