module blink_top (
	input clk_50,
	input reset_btn,
	output [3:0] led
	);
	
	
	
nios_old nios_instance (
		.clk_clk (clk_50),       //   clk.clk
		.gpio_export (led),   //  gpio.export
		.reset_reset_n (reset_btn) // reset.reset_n
	);

endmodule